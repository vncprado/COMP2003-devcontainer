module and_gate (
    output logic y,
    input logic a, b
);
    
endmodule